----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:22:45 04/22/2009 
-- Design Name: 
-- Module Name:    mux2_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity mux2_1 is
	port(I0, I1, S : in STD_LOGIC;
	     o : out STD_LOGIC);
end mux2_1;

architecture multiplexer of mux2_1 is
begin
	sel: process (S, I0, I1) 
	begin
		if (S = '0') then
			o <= I0;
		else
			o <= I1;
		end if;
	end process;
	SCLK_pull: PULLDOWN port map(O=>o);
end multiplexer;

